library verilog;
use verilog.vl_types.all;
entity lab9part1_vlg_vec_tst is
end lab9part1_vlg_vec_tst;
