library verilog;
use verilog.vl_types.all;
entity lab11part1_vlg_vec_tst is
end lab11part1_vlg_vec_tst;
