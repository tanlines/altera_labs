library verilog;
use verilog.vl_types.all;
entity part4_vlg_vec_tst is
end part4_vlg_vec_tst;
