library verilog;
use verilog.vl_types.all;
entity part1_vlg_vec_tst is
end part1_vlg_vec_tst;
