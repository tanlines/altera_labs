library verilog;
use verilog.vl_types.all;
entity part2_vlg_vec_tst is
end part2_vlg_vec_tst;
