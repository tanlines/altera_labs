library verilog;
use verilog.vl_types.all;
entity countertest_vlg_vec_tst is
end countertest_vlg_vec_tst;
