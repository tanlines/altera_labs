library verilog;
use verilog.vl_types.all;
entity part4_vlg_check_tst is
    port(
        Q_a             : in     vl_logic;
        Q_b             : in     vl_logic;
        Q_c             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end part4_vlg_check_tst;
